library verilog;
use verilog.vl_types.all;
entity EDA2_tb is
end EDA2_tb;
